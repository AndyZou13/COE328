library verilog;
use verilog.vl_types.all;
entity john_vlg_vec_tst is
end john_vlg_vec_tst;
