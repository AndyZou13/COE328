library verilog;
use verilog.vl_types.all;
entity seg7_vlg_vec_tst is
end seg7_vlg_vec_tst;
